��  CCircuit��  CSerializeHack           ��  CPart              ��� 	 CLogicOut�� 	 CTerminal  ����              @            ����          ��    �
�  ��               �            ��            ��    ��  CLogicIn�� 	 CLatchKey  � �� �         
�  � �� �                            � �� �         ����     ��  � 	�          
�  � �                             � �          ����     ��  CNOR
�  � ��               �          
�  � ��                          
�  �1�              @            ��           ��    �
�  �                           
�  �  !              @          
�  1               �            $           ��                  ���  CWire  X�       �  0Y       ��� 
 CCrossOver  VL\T        XYy        �$�  VL\T        � PiQ       �  � xYy       �  � x� �        �  � �� �       �  h���       �  0�i�       �  hPi�        �  �  � Q        �  �  � !       �  � �� �       �  � �                     �                             +   !    0   1  *   0    ,  1   /    " "   # # ' ! ( & % . - ) # ( * )  ,   - & + / & .                  �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 