��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  �)7    EX-NOR      �  ���    EX-OR      �  �!/    NOR      �  � �� �    NOT      �  � 9� G    NAND      �  � �� �    OR      �  � )� 7    AND          �   �     ��� 	 CLogicOut�� 	 CTerminal  �p�q               �            �h�x           ��    ��  CLogicIn�� 	 CLatchKey  �y��         �  ����                            �|��         ����     ��  CAND�  8�M�              @          �  8�M�                          �  d�y�               �            L�d�           ��    ��  COR�  �h�i               �          �  �x�y               �          �  �p�q               �            �d�|            ��    ��  �I�W     #   �  �P�Q              @            �L�T     %   ����     ��  8PMQ               �          �  8`Ma              @          �  dXyY               �            LLdd     '      ��    �� 	 CInverter�  ����                          �  �!�              @            �t�     ,      ��    *��  �P�Q              @          �  P!Q               �            �D\     /      ��    ��   �5�              @            4�D�     2     ��    ��  ����      3   �  ����                            ����     5    ����     ��  ����     6   �  ����              @            ����     8   ����     ��  CXOR�  ����              @          �  ����                          �  ��              @            ���     ;      ��    ��   P5Q               �            4HDX     ?      ��    ��  �Y�g     @   �  �`�a              @            �\�d     B   ����     ��  �9�G      C   �  �@�A                            �<�D     E    ����     ��  CNOR�  �H�I                          �  �X�Y              @          �  PQ               �            �D\     H      ��    ��  �-�     
          �            ,�<�     L      ��    ��  � �� �     M   �  � �� �              @            � �� �     O   ����     *��  � �� �              @          �  � ��     
          �            � �� �     Q      ��    ��  h-i               �            ,`<p     T      ��    ��  � y� �     U   �  � �� �     	         @            � |� �     W   ����     ��  � I� W     X   �  � P� Q              @            � L� T     Z   ����     ��  CNAND�  � `� a              @          �  � p� q     	         @          �  � hi               �            � \� t     ]      ��    ��  �%�              @            $�4�     a     ��    ��  � �      b   �  � � 	              @            � �      d   ����     ��  � �� �      e   �  � �� �                            � �� �     g    ����     ��  � �� �                          �  � �� �              @          �  � �	�              @            � �� �     i      ��    ��  XY              @            P,`     m     ��    ��  � i� w     n   �  � p� q              @            � l� t     p   ����     ��  � P� Q              @          �  � `� a              @          �  � XY              @            � L� d     r      ��    ��  � 9� G     u   �  � @� A              @            � <� D     w   ����         �   �     ���  CWire  �p�q      y�  ��9�      y��� 
 CCrossOver  ����        ����       y�}�  ����        ��9�      y�  �P�i       y�  �h�i      y�  �h��       y�  ����      y�  �x��       y�  x���      y�  �X�i       y�  xX�Y      y�  �P�Q      y�   �9�      y�  8`9�       y�   P9Q      y�  �!�      y�  ����       y�  ����      y�  ����       y�  ����      y�  P!Q      y�  �X�a       y�  �`�a      y�  �@�I       y�  �@�A      y�  ��     
 y�  � �� �       y�  � �� �      y�  hi      y�  � p� �      	 y�  � �� �     	 y�  � P� a       y�  � P� Q      y�  ��      y�  � �� �       y�  � �� �      y�  � �� 	       y�  � � 	      y�   X	Y      y�  � `� q       y�  � p� q      y�  � @� Q       y�  � @� A          �   �     �    �   �         �   �      z    �     {    �   �   ! � ! " " z % % � ' � ' ( � ( ) ) � , � , - - � / � / 0 0 � 2 � 2 5 5 � 8 8 � ; � ; < � < = = � ? � ? B B � E E � H � H I � I J J � L � L O O � Q � Q R R � T � T W W � Z Z � ] � ] ^ � ^ _ _ � a � a d d � g g � i � i j � j k k � m � m p p � r � r s � s t t � w w � "  |  | �  {  ~ �  % � � � �  | , ! �  � �   ) � � / - � ( � 0 ' = 2 < � 5 � � ; 8 � J ? I � B � � H E � R L Q � O � _ T ^ � W � � ] Z � k a � i g � j � d � t m s � p � � r w �             �$s�        @!Muhammad Rifqi Athallah 202031234    +        @            @    "V  (      ��                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 