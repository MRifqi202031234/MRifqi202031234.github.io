��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  ��    Output      �  �)�7    A      �  �9�G    B      �  �I�W    A      �  �Y�g    B      �  q)|7    A      �  q9|G    B      �  qI|W    A      �  qY|g    B      �  IYSg    1      �  IISW    1      �  I9SG    0      �  � �� �    C      �  � �� �    B      �  � y� �    A      �  ����    Output      �  I)S7    0      �  q|    B      �  IT    A      �  ��    Output      �  � )� 7    B      �  � 	�     A                  ���  CAND�� 	 CTerminal  x���               �          !�  x���                          !�  ����     	          �            ����     "      ��    �� 	 CLogicOut!�  ����     	          �            ����     '      ��    ��  CLogicIn�� 	 CLatchKey  � �� �      )   !�  ��                            � ��     ,    ����     (�*�  � �� �      -   !�  ��                            � ��     /    ����     (�*�  � y� �      0   !�  ��                            � |�     2    ����     �!�  (�=�                          !�  (�=�                          !�  T�i�               �            <�T�     4      ��    %�!�  p �!              @            ��(     8     ��    (�*�  � )� 7     9   !�  01              @            � ,4     ;   ����     (�*�  � 	�      <   !�                @            �      >   ����     �!�  (=              @          !�  ((=)              @          !�  T i!              @            <T,     @      ��                ���  CWire  ����      	 D�  ����     	 D�  �y�      D�  h�y�      D�  h�i�       D�  (�)�       D�  �)�      D�  (�)�       D�  �)�      D�  )      D�  h q!      D�  (()1       D�  0)1      D�  ()                   �                        " H " # G # $ $ F ' E ' , , G / / K 2 2 M 4 L 4 5 J 5 6 6 I 8 O 8 ; ; Q > > N @ R @ A P A B B O ' F $ E , # I " 6 H 5 K / J M 4 2 L > R B 8 A Q ; P N @             �$s�        @Praktikum 4    +        @            @    "V  (      �8                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 